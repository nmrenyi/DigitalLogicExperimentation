library verilog;
use verilog.vl_types.all;
entity CarryLookAheadAdder_vlg_vec_tst is
end CarryLookAheadAdder_vlg_vec_tst;
