library verilog;
use verilog.vl_types.all;
entity TEF_vlg_vec_tst is
end TEF_vlg_vec_tst;
