library verilog;
use verilog.vl_types.all;
entity Counter_vlg_vec_tst is
end Counter_vlg_vec_tst;
