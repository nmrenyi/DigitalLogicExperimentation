library verilog;
use verilog.vl_types.all;
entity Light_vlg_vec_tst is
end Light_vlg_vec_tst;
