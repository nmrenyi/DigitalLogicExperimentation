library verilog;
use verilog.vl_types.all;
entity DigitalLife_vlg_vec_tst is
end DigitalLife_vlg_vec_tst;
