library verilog;
use verilog.vl_types.all;
entity Serial4FullAdder_vlg_vec_tst is
end Serial4FullAdder_vlg_vec_tst;
